CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 9
0 71 1920 939
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
36 C:\Program Files (x86)\CM60S\BOM.DAT
0 7
0 71 1920 939
144179218 0
0
6 Title:
5 Name:
0
0
0
19
11 Multimeter~
205 480 186 0 21 21
0 11 12 13 9 0 0 0 0 0
32 57 57 50 46 50 117 65 0 0
0 86
0
0 0 16464 0
6 1.000u
-21 -19 21 -11
3 MM0
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
7 Ground~
168 771 446 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
13 Var Resistor~
219 876 240 0 3 7
0 3 4 14
0
0 0 848 90
7 10k 20%
10 -5 59 3
3 POT
24 -14 45 -6
0
0
30 %DA %1 %2 2000
%DB %2 %3 8000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 512 1 0 0 0
1 R
3618 0 0
0
0
7 Ground~
168 1019 311 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
11 Multimeter~
205 979 257 0 21 21
0 3 15 16 2 0 0 0 0 0
32 53 46 48 48 48 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
7 Ground~
168 425 323 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
9 V Source~
197 425 264 0 2 5
0 11 2
0
0 0 17264 0
2 9V
17 0 31 8
3 Vs1
13 -10 34 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
2 Vs
9914 0 0
0
0
8 Op-Amp5~
219 814 338 0 5 11
0 6 5 9 2 3
0
0 0 848 0
5 LM358
15 -25 50 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 1216257740
88 0 0 256 2 1 1 0
1 U
3747 0 0
0
0
7 Ground~
168 831 389 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 647 445 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
7 Ground~
168 525 446 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
9 Resistor~
219 771 390 0 3 5
0 2 6 -1
0
0 0 880 90
4 100k
2 -1 30 7
2 R7
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 820 238 0 2 5
0 5 4
0
0 0 880 0
4 132k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 718 344 0 2 5
0 7 6
0
0 0 880 0
4 100k
-13 18 15 26
2 R5
-7 6 7 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
9 Resistor~
219 706 332 0 2 5
0 8 5
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 647 390 0 3 5
0 2 7 -1
0
0 0 880 90
3 20k
5 0 26 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 525 387 0 3 5
0 2 8 -1
0
0 0 880 90
2 22
10 -1 24 7
3 LDR
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 647 268 0 2 5
0 7 9
0
0 0 880 90
3 20k
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 526 270 0 2 5
0 8 9
0
0 0 880 90
3 20k
5 0 26 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
22
4 1 2 0 0 4096 0 5 4 0 0 4
1004 280
1004 297
1019 297
1019 305
1 1 2 0 0 4096 0 2 12 0 0 2
771 440
771 408
1 0 3 0 0 4096 0 3 0 0 5 2
880 254
880 296
2 2 4 0 0 4224 0 3 13 0 0 2
868 238
838 238
1 5 3 0 0 8320 0 5 8 0 0 5
954 280
954 296
880 296
880 338
832 338
1 2 2 0 0 0 0 6 7 0 0 2
425 317
425 285
0 1 5 0 0 4224 0 0 13 16 0 3
756 332
756 238
802 238
2 0 6 0 0 4096 0 12 0 0 15 2
771 372
771 344
1 0 7 0 0 4096 0 14 0 0 19 2
700 344
647 344
1 0 8 0 0 20608 0 15 0 0 20 6
688 332
657 332
657 325
637 325
637 332
525 332
4 2 9 0 0 24576 0 1 19 0 0 7
505 209
504 209
504 209
527 209
527 209
526 209
526 252
1 4 2 0 0 0 0 9 8 0 0 4
831 383
831 366
814 366
814 351
0 3 9 0 0 32768 0 0 8 17 0 10
647 209
685 209
685 260
747 260
747 251
768 251
768 260
815 260
815 325
814 325
0 0 10 0 0 0 0 0 0 0 0 2
909 238
909 238
2 1 6 0 0 4224 0 14 8 0 0 2
736 344
796 344
2 2 5 0 0 0 0 15 8 0 0 2
724 332
796 332
2 0 9 0 0 8320 0 18 0 0 11 3
647 250
647 209
527 209
1 1 11 0 0 4224 0 7 1 0 0 3
425 243
425 209
455 209
1 2 7 0 0 4224 0 18 16 0 0 2
647 286
647 372
1 2 8 0 0 0 0 19 17 0 0 3
526 288
525 288
525 369
1 1 2 0 0 0 0 10 16 0 0 2
647 439
647 408
1 1 2 0 0 4224 0 11 17 0 0 2
525 440
525 405
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
17367698 1210432 100 100 0 0
0 0 0 0
0 71 161 141
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 5
0
33947850 8534080 100 100 0 0
77 66 1877 396
0 555 1920 1039
1877 66
77 66
1877 66
1877 396
0 0
5e-006 0 5e-006 0 5e-006 5e-006
12393 0
4 1e-006 5
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
